1��ش ��1���� �� � ~��1���� �� � ���� ~  �3                                                                                                                                                                                                                                                                                                                                                                                                                                                                         U��9`1������&�� �  &�� �Z�&�� �  &�� ���&�� �  &�� �H�&�� �  &�� �8�&�� �  &�� ��&�� �  &�� ��&�� �  &�� ��&�� �  &�� ��&�� �  &�� �&�� �  &�� ��~&�� �  &�� ���&�� �  &�� �ـ&�� �  &�� a�`�)�.�����1����6����� ������  ��.t�Ί< t���!�#��B��a�`� �*��)S�.�����1����6����� ���[���  ��.t"�Ί< t��Q�,��ƹ	 �Y�0	�t��B�ٸŅ�!�#� �ˀ��t,�˃�	� ��)�.�����1����6������G�������NS�*�1���+��[�ˊW	� �ӈ*�����!����"�?nt!�?yu�u��5��@ �u��\C�߾,��	 �a�Q�%��P���%X9�t �Ɖ��t� ��  Y�`� ��a�RQSP�߻
 1�1���RA�� u�X0���0��X[YZ�P�ƹ  ��tA��X�`�ǹ  � �9�tA��a�`�߹  ��t%� �<u�� t��<t<t�A��I9�t�O�ִ��� ���
�a�`�����
�a�`�Ƭ�t����a�`��1���S1۹��S� � �a�`1���r2� ���&�ػ �!��/�� ���&�ػ �!��/����&�ػ �!a�`R1ҋ����BR1ҋ�������XZ���������a����1��؎��2�'�<��)��!�u��\�����)��!����*��!�u��*��!����)��!����"�? tӻ������0�� �� �������0�� ta�������0�� t8�������0�� t]�������0�� �� �����0�� tY�������0�� t#��#�*�� ��2�#�b��#����1�#�V��'�Q��3�#�ꅻ)��!�#�@��#�4�#�7��#����)��!�#�(��*�<t�5��u��@ �+�1���*�����#����)��!�#����#����!�u��!�#������� �$�1�����?������6���        A: > \ Directory does not have a parent directory! Already at root directory! This is a directory!
Would you like to change your current working directory? [y/n]:  MonsterOS Version 1.1
Copyright (C) 2014 Daniel Lopez. Licensed Under The Simplified BSD License
 
MonsterOS  Welcome to the MonsterOS shell prompt.

MonsterOS shell prompt contains only two internal commands: help, clear, and list.
This means that MonsterOS treats everything else that is not the help/clear command as an external command.
An external command is basically a filename of a file stored on the disk.
If the file is located on the disk it is executed if it is a program; else it is treated a text file and its contents are displayed.
If no file is found then a error message is displayed. help clear list poweroff date pwd .. Invalid Internal / External Command! Machine failed to shutdown!!!
Error: APM May Not Be Supported                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �System16 ver.com  	dbug.com 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               krnl.sys                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ���� ��!�MonsterOS Version 1.1                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 RQSP�;��!X�^��&�^��!��	��@��!X�^��&�^��!�� ��E��!X�^��&�^��!�� ��J��!X�^��&�^��!�� ��O��!X�^��&�^��!�� ��T��!X�^��&�^��!�� ��Y��!X�^��&�^��!�� ��AX:  BX:  CX:  DX:  CS:  DS:  ES:                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �#����!�#�Error: This is a system file! Cannot be executed!                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     